module top(
    input [1:0] sel,
    input [17:0] DIA, DIB,
    output [17:0] DOA, DOB,
    input [13:0] ADA, ADB,
    input CEA, OCEA, CLKA, WEA, CSA2, CSA1, CSA0, RSTA,
    input CEB, OCEB, CLKB, WEB, CSB2, CSB1, CSB0, RSTB
);

wire [17:0] DOA_I[0:2];
wire [17:0] DOB_I[0:2];

DP8KC  #(
    .WRITEMODE_A("NORMAL"), .WRITEMODE_B("NORMAL")
) ebr_NORMAL_NORMAL (
    .DIA0(DIA[0]), .DIA1(DIA[1]), .DIA2(DIA[2]), .DIA3(DIA[3]), .DIA4(DIA[4]), .DIA5(DIA[5]), .DIA6(DIA[6]), .DIA7(DIA[7]), .DIA8(DIA[8]),
    .DIB0(DIB[0]), .DIB1(DIB[1]), .DIB2(DIB[2]), .DIB3(DIB[3]), .DIB4(DIB[4]), .DIB5(DIB[5]), .DIB6(DIB[6]), .DIB7(DIB[7]), .DIB8(DIB[8]),
    .ADA0(ADA[0]), .ADA1(ADA[1]), .ADA2(ADA[2]), .ADA3(ADA[3]), .ADA4(ADA[4]), .ADA5(ADA[5]), .ADA6(ADA[6]), .ADA7(ADA[7]), .ADA8(ADA[8]), .ADA9(ADA[9]), .ADA10(ADA[10]), .ADA11(ADA[11]), .ADA12(ADA[12]),
    .ADB0(ADB[0]), .ADB1(ADB[1]), .ADB2(ADB[2]), .ADB3(ADB[3]), .ADB4(ADB[4]), .ADB5(ADB[5]), .ADB6(ADB[6]), .ADB7(ADB[7]), .ADB8(ADB[8]), .ADB9(ADB[9]), .ADB10(ADB[10]), .ADB11(ADB[11]), .ADB12(ADB[12]),
    .DOA0(DOA_I[0][0]), .DOA1(DOA_I[0][1]), .DOA2(DOA_I[0][2]), .DOA3(DOA_I[0][3]), .DOA4(DOA_I[0][4]), .DOA5(DOA_I[0][5]), .DOA6(DOA_I[0][6]), .DOA7(DOA_I[0][7]), .DOA8(DOA_I[0][8]),
    .DOB0(DOB_I[0][0]), .DOB1(DOB_I[0][1]), .DOB2(DOB_I[0][2]), .DOB3(DOB_I[0][3]), .DOB4(DOB_I[0][4]), .DOB5(DOB_I[0][5]), .DOB6(DOB_I[0][6]), .DOB7(DOB_I[0][7]), .DOB8(DOB_I[0][8]),
    .CEA(CEA), .OCEA(OCEA), .CLKA(CLKA), .WEA(WEA), .CSA2(CSA2), .CSA1(CSA1), .CSA0(CSA0), .RSTA(RSTA),
    .CEB(CEB), .OCEB(OCEB), .CLKB(CLKB), .WEB(WEB), .CSB2(CSB2), .CSB1(CSB1), .CSB0(CSB0), .RSTB(RSTB)
);

DP8KC  #(
    .WRITEMODE_A("NORMAL"), .WRITEMODE_B("READBEFOREWRITE")
) ebr_NORMAL_READBEFOREWRITE (
    .DIA0(DIA[0]), .DIA1(DIA[1]), .DIA2(DIA[2]), .DIA3(DIA[3]), .DIA4(DIA[4]), .DIA5(DIA[5]), .DIA6(DIA[6]), .DIA7(DIA[7]), .DIA8(DIA[8]),
    .DIB0(DIB[0]), .DIB1(DIB[1]), .DIB2(DIB[2]), .DIB3(DIB[3]), .DIB4(DIB[4]), .DIB5(DIB[5]), .DIB6(DIB[6]), .DIB7(DIB[7]), .DIB8(DIB[8]),
    .ADA0(ADA[0]), .ADA1(ADA[1]), .ADA2(ADA[2]), .ADA3(ADA[3]), .ADA4(ADA[4]), .ADA5(ADA[5]), .ADA6(ADA[6]), .ADA7(ADA[7]), .ADA8(ADA[8]), .ADA9(ADA[9]), .ADA10(ADA[10]), .ADA11(ADA[11]), .ADA12(ADA[12]),
    .ADB0(ADB[0]), .ADB1(ADB[1]), .ADB2(ADB[2]), .ADB3(ADB[3]), .ADB4(ADB[4]), .ADB5(ADB[5]), .ADB6(ADB[6]), .ADB7(ADB[7]), .ADB8(ADB[8]), .ADB9(ADB[9]), .ADB10(ADB[10]), .ADB11(ADB[11]), .ADB12(ADB[12]),
    .DOA0(DOA_I[1][0]), .DOA1(DOA_I[1][1]), .DOA2(DOA_I[1][2]), .DOA3(DOA_I[1][3]), .DOA4(DOA_I[1][4]), .DOA5(DOA_I[1][5]), .DOA6(DOA_I[1][6]), .DOA7(DOA_I[1][7]), .DOA8(DOA_I[1][8]),
    .DOB0(DOB_I[1][0]), .DOB1(DOB_I[1][1]), .DOB2(DOB_I[1][2]), .DOB3(DOB_I[1][3]), .DOB4(DOB_I[1][4]), .DOB5(DOB_I[1][5]), .DOB6(DOB_I[1][6]), .DOB7(DOB_I[1][7]), .DOB8(DOB_I[1][8]),
    .CEA(CEA), .OCEA(OCEA), .CLKA(CLKA), .WEA(WEA), .CSA2(CSA2), .CSA1(CSA1), .CSA0(CSA0), .RSTA(RSTA),
    .CEB(CEB), .OCEB(OCEB), .CLKB(CLKB), .WEB(WEB), .CSB2(CSB2), .CSB1(CSB1), .CSB0(CSB0), .RSTB(RSTB)
);

DP8KC  #(
   .WRITEMODE_A("NORMAL"), .WRITEMODE_B("WRITETHROUGH")
) ebr_NORMAL_WRITETHROUGH (
    .DIA0(DIA[0]), .DIA1(DIA[1]), .DIA2(DIA[2]), .DIA3(DIA[3]), .DIA4(DIA[4]), .DIA5(DIA[5]), .DIA6(DIA[6]), .DIA7(DIA[7]), .DIA8(DIA[8]),
    .DIB0(DIB[0]), .DIB1(DIB[1]), .DIB2(DIB[2]), .DIB3(DIB[3]), .DIB4(DIB[4]), .DIB5(DIB[5]), .DIB6(DIB[6]), .DIB7(DIB[7]), .DIB8(DIB[8]),
    .ADA0(ADA[0]), .ADA1(ADA[1]), .ADA2(ADA[2]), .ADA3(ADA[3]), .ADA4(ADA[4]), .ADA5(ADA[5]), .ADA6(ADA[6]), .ADA7(ADA[7]), .ADA8(ADA[8]), .ADA9(ADA[9]), .ADA10(ADA[10]), .ADA11(ADA[11]), .ADA12(ADA[12]),
    .ADB0(ADB[0]), .ADB1(ADB[1]), .ADB2(ADB[2]), .ADB3(ADB[3]), .ADB4(ADB[4]), .ADB5(ADB[5]), .ADB6(ADB[6]), .ADB7(ADB[7]), .ADB8(ADB[8]), .ADB9(ADB[9]), .ADB10(ADB[10]), .ADB11(ADB[11]), .ADB12(ADB[12]),
    .DOA0(DOA_I[2][0]), .DOA1(DOA_I[2][1]), .DOA2(DOA_I[2][2]), .DOA3(DOA_I[2][3]), .DOA4(DOA_I[2][4]), .DOA5(DOA_I[2][5]), .DOA6(DOA_I[2][6]), .DOA7(DOA_I[2][7]), .DOA8(DOA_I[2][8]),
    .DOB0(DOB_I[2][0]), .DOB1(DOB_I[2][1]), .DOB2(DOB_I[2][2]), .DOB3(DOB_I[2][3]), .DOB4(DOB_I[2][4]), .DOB5(DOB_I[2][5]), .DOB6(DOB_I[2][6]), .DOB7(DOB_I[2][7]), .DOB8(DOB_I[2][8]),
    .CEA(CEA), .OCEA(OCEA), .CLKA(CLKA), .WEA(WEA), .CSA2(CSA2), .CSA1(CSA1), .CSA0(CSA0), .RSTA(RSTA),
    .CEB(CEB), .OCEB(OCEB), .CLKB(CLKB), .WEB(WEB), .CSB2(CSB2), .CSB1(CSB1), .CSB0(CSB0), .RSTB(RSTB)
);




assign DOA = DOA_I[sel];
assign DOB = DOB_I[sel];


endmodule
