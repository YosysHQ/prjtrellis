module ILVDS(input A, AN, output Z);
    assign Z = A; //yeah, they really did this, no checking of AN
endmodule // ILVDS

    
