module top(output f);
    assign f = 0;
endmodule
