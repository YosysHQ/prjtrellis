module top(
    input [1:0] sel,
    input [17:0] DIA, DIB,
    output [17:0] DOA, DOB,
    input [13:0] ADA, ADB,
    input CEA, OCEA, CLKA, WEA, CSA2, CSA1, CSA0, RSTA,
    input CEB, OCEB, CLKB, WEB, CSB2, CSB1, CSB0, RSTB
);

wire [17:0] DOA_I[0:3];
wire [17:0] DOB_I[0:3];

DP16KD  #(
    .REGMODE_A("NOREG"), .REGMODE_B("NOREG")
) ebr_NOREG_NOREG (
    .DIA0(DIA[0]), .DIA1(DIA[1]), .DIA2(DIA[2]), .DIA3(DIA[3]), .DIA4(DIA[4]), .DIA5(DIA[5]), .DIA6(DIA[6]), .DIA7(DIA[7]), .DIA8(DIA[8]), .DIA9(DIA[9]), .DIA10(DIA[10]), .DIA11(DIA[11]), .DIA12(DIA[12]), .DIA13(DIA[13]), .DIA14(DIA[14]), .DIA15(DIA[15]), .DIA16(DIA[16]), .DIA17(DIA[17]),
    .DIB0(DIB[0]), .DIB1(DIB[1]), .DIB2(DIB[2]), .DIB3(DIB[3]), .DIB4(DIB[4]), .DIB5(DIB[5]), .DIB6(DIB[6]), .DIB7(DIB[7]), .DIB8(DIB[8]), .DIB9(DIB[9]), .DIB10(DIB[10]), .DIB11(DIB[11]), .DIB12(DIB[12]), .DIB13(DIB[13]), .DIB14(DIB[14]), .DIB15(DIB[15]), .DIB16(DIB[16]), .DIB17(DIB[17]),
    .ADA0(ADA[0]), .ADA1(ADA[1]), .ADA2(ADA[2]), .ADA3(ADA[3]), .ADA4(ADA[4]), .ADA5(ADA[5]), .ADA6(ADA[6]), .ADA7(ADA[7]), .ADA8(ADA[8]), .ADA9(ADA[9]), .ADA10(ADA[10]), .ADA11(ADA[11]), .ADA12(ADA[12]), .ADA13(ADA[13]),
    .ADB0(ADB[0]), .ADB1(ADB[1]), .ADB2(ADB[2]), .ADB3(ADB[3]), .ADB4(ADB[4]), .ADB5(ADB[5]), .ADB6(ADB[6]), .ADB7(ADB[7]), .ADB8(ADB[8]), .ADB9(ADB[9]), .ADB10(ADB[10]), .ADB11(ADB[11]), .ADB12(ADB[12]), .ADB13(ADB[13]),
    .DOA0(DOA_I[0][0]), .DOA1(DOA_I[0][1]), .DOA2(DOA_I[0][2]), .DOA3(DOA_I[0][3]), .DOA4(DOA_I[0][4]), .DOA5(DOA_I[0][5]), .DOA6(DOA_I[0][6]), .DOA7(DOA_I[0][7]), .DOA8(DOA_I[0][8]), .DOA9(DOA_I[0][9]), .DOA10(DOA_I[0][10]), .DOA11(DOA_I[0][11]), .DOA12(DOA_I[0][12]), .DOA13(DOA_I[0][13]), .DOA14(DOA_I[0][14]), .DOA15(DOA_I[0][15]), .DOA16(DOA_I[0][16]), .DOA17(DOA_I[0][17]),
    .DOB0(DOB_I[0][0]), .DOB1(DOB_I[0][1]), .DOB2(DOB_I[0][2]), .DOB3(DOB_I[0][3]), .DOB4(DOB_I[0][4]), .DOB5(DOB_I[0][5]), .DOB6(DOB_I[0][6]), .DOB7(DOB_I[0][7]), .DOB8(DOB_I[0][8]), .DOB9(DOB_I[0][9]), .DOB10(DOB_I[0][10]), .DOB11(DOB_I[0][11]), .DOB12(DOB_I[0][12]), .DOB13(DOB_I[0][13]), .DOB14(DOB_I[0][14]), .DOB15(DOB_I[0][15]), .DOB16(DOB_I[0][16]), .DOB17(DOB_I[0][17]),
    .CEA(CEA), .OCEA(OCEA), .CLKA(CLKA), .WEA(WEA), .CSA2(CSA2), .CSA1(CSA1), .CSA0(CSA0), .RSTA(RSTA),
    .CEB(CEB), .OCEB(OCEB), .CLKB(CLKB), .WEB(WEB), .CSB2(CSB2), .CSB1(CSB1), .CSB0(CSB0), .RSTB(RSTB)
);

DP16KD  #(
    .REGMODE_A("NOREG"), .REGMODE_B("OUTREG")
) ebr_NOREG_OUTREG (
    .DIA0(DIA[0]), .DIA1(DIA[1]), .DIA2(DIA[2]), .DIA3(DIA[3]), .DIA4(DIA[4]), .DIA5(DIA[5]), .DIA6(DIA[6]), .DIA7(DIA[7]), .DIA8(DIA[8]), .DIA9(DIA[9]), .DIA10(DIA[10]), .DIA11(DIA[11]), .DIA12(DIA[12]), .DIA13(DIA[13]), .DIA14(DIA[14]), .DIA15(DIA[15]), .DIA16(DIA[16]), .DIA17(DIA[17]),
    .DIB0(DIB[0]), .DIB1(DIB[1]), .DIB2(DIB[2]), .DIB3(DIB[3]), .DIB4(DIB[4]), .DIB5(DIB[5]), .DIB6(DIB[6]), .DIB7(DIB[7]), .DIB8(DIB[8]), .DIB9(DIB[9]), .DIB10(DIB[10]), .DIB11(DIB[11]), .DIB12(DIB[12]), .DIB13(DIB[13]), .DIB14(DIB[14]), .DIB15(DIB[15]), .DIB16(DIB[16]), .DIB17(DIB[17]),
    .ADA0(ADA[0]), .ADA1(ADA[1]), .ADA2(ADA[2]), .ADA3(ADA[3]), .ADA4(ADA[4]), .ADA5(ADA[5]), .ADA6(ADA[6]), .ADA7(ADA[7]), .ADA8(ADA[8]), .ADA9(ADA[9]), .ADA10(ADA[10]), .ADA11(ADA[11]), .ADA12(ADA[12]), .ADA13(ADA[13]),
    .ADB0(ADB[0]), .ADB1(ADB[1]), .ADB2(ADB[2]), .ADB3(ADB[3]), .ADB4(ADB[4]), .ADB5(ADB[5]), .ADB6(ADB[6]), .ADB7(ADB[7]), .ADB8(ADB[8]), .ADB9(ADB[9]), .ADB10(ADB[10]), .ADB11(ADB[11]), .ADB12(ADB[12]), .ADB13(ADB[13]),
    .DOA0(DOA_I[1][0]), .DOA1(DOA_I[1][1]), .DOA2(DOA_I[1][2]), .DOA3(DOA_I[1][3]), .DOA4(DOA_I[1][4]), .DOA5(DOA_I[1][5]), .DOA6(DOA_I[1][6]), .DOA7(DOA_I[1][7]), .DOA8(DOA_I[1][8]), .DOA9(DOA_I[1][9]), .DOA10(DOA_I[1][10]), .DOA11(DOA_I[1][11]), .DOA12(DOA_I[1][12]), .DOA13(DOA_I[1][13]), .DOA14(DOA_I[1][14]), .DOA15(DOA_I[1][15]), .DOA16(DOA_I[1][16]), .DOA17(DOA_I[1][17]),
    .DOB0(DOB_I[1][0]), .DOB1(DOB_I[1][1]), .DOB2(DOB_I[1][2]), .DOB3(DOB_I[1][3]), .DOB4(DOB_I[1][4]), .DOB5(DOB_I[1][5]), .DOB6(DOB_I[1][6]), .DOB7(DOB_I[1][7]), .DOB8(DOB_I[1][8]), .DOB9(DOB_I[1][9]), .DOB10(DOB_I[1][10]), .DOB11(DOB_I[1][11]), .DOB12(DOB_I[1][12]), .DOB13(DOB_I[1][13]), .DOB14(DOB_I[1][14]), .DOB15(DOB_I[1][15]), .DOB16(DOB_I[1][16]), .DOB17(DOB_I[1][17]),
    .CEA(CEA), .OCEA(OCEA), .CLKA(CLKA), .WEA(WEA), .CSA2(CSA2), .CSA1(CSA1), .CSA0(CSA0), .RSTA(RSTA),
    .CEB(CEB), .OCEB(OCEB), .CLKB(CLKB), .WEB(WEB), .CSB2(CSB2), .CSB1(CSB1), .CSB0(CSB0), .RSTB(RSTB)
);

DP16KD  #(
    .REGMODE_A("OUTREG"), .REGMODE_B("NOREG")
) ebr_OUTREG_NOREG (
    .DIA0(DIA[0]), .DIA1(DIA[1]), .DIA2(DIA[2]), .DIA3(DIA[3]), .DIA4(DIA[4]), .DIA5(DIA[5]), .DIA6(DIA[6]), .DIA7(DIA[7]), .DIA8(DIA[8]), .DIA9(DIA[9]), .DIA10(DIA[10]), .DIA11(DIA[11]), .DIA12(DIA[12]), .DIA13(DIA[13]), .DIA14(DIA[14]), .DIA15(DIA[15]), .DIA16(DIA[16]), .DIA17(DIA[17]),
    .DIB0(DIB[0]), .DIB1(DIB[1]), .DIB2(DIB[2]), .DIB3(DIB[3]), .DIB4(DIB[4]), .DIB5(DIB[5]), .DIB6(DIB[6]), .DIB7(DIB[7]), .DIB8(DIB[8]), .DIB9(DIB[9]), .DIB10(DIB[10]), .DIB11(DIB[11]), .DIB12(DIB[12]), .DIB13(DIB[13]), .DIB14(DIB[14]), .DIB15(DIB[15]), .DIB16(DIB[16]), .DIB17(DIB[17]),
    .ADA0(ADA[0]), .ADA1(ADA[1]), .ADA2(ADA[2]), .ADA3(ADA[3]), .ADA4(ADA[4]), .ADA5(ADA[5]), .ADA6(ADA[6]), .ADA7(ADA[7]), .ADA8(ADA[8]), .ADA9(ADA[9]), .ADA10(ADA[10]), .ADA11(ADA[11]), .ADA12(ADA[12]), .ADA13(ADA[13]),
    .ADB0(ADB[0]), .ADB1(ADB[1]), .ADB2(ADB[2]), .ADB3(ADB[3]), .ADB4(ADB[4]), .ADB5(ADB[5]), .ADB6(ADB[6]), .ADB7(ADB[7]), .ADB8(ADB[8]), .ADB9(ADB[9]), .ADB10(ADB[10]), .ADB11(ADB[11]), .ADB12(ADB[12]), .ADB13(ADB[13]),
    .DOA0(DOA_I[2][0]), .DOA1(DOA_I[2][1]), .DOA2(DOA_I[2][2]), .DOA3(DOA_I[2][3]), .DOA4(DOA_I[2][4]), .DOA5(DOA_I[2][5]), .DOA6(DOA_I[2][6]), .DOA7(DOA_I[2][7]), .DOA8(DOA_I[2][8]), .DOA9(DOA_I[2][9]), .DOA10(DOA_I[2][10]), .DOA11(DOA_I[2][11]), .DOA12(DOA_I[2][12]), .DOA13(DOA_I[2][13]), .DOA14(DOA_I[2][14]), .DOA15(DOA_I[2][15]), .DOA16(DOA_I[2][16]), .DOA17(DOA_I[2][17]),
    .DOB0(DOB_I[2][0]), .DOB1(DOB_I[2][1]), .DOB2(DOB_I[2][2]), .DOB3(DOB_I[2][3]), .DOB4(DOB_I[2][4]), .DOB5(DOB_I[2][5]), .DOB6(DOB_I[2][6]), .DOB7(DOB_I[2][7]), .DOB8(DOB_I[2][8]), .DOB9(DOB_I[2][9]), .DOB10(DOB_I[2][10]), .DOB11(DOB_I[2][11]), .DOB12(DOB_I[2][12]), .DOB13(DOB_I[2][13]), .DOB14(DOB_I[2][14]), .DOB15(DOB_I[2][15]), .DOB16(DOB_I[2][16]), .DOB17(DOB_I[2][17]),
    .CEA(CEA), .OCEA(OCEA), .CLKA(CLKA), .WEA(WEA), .CSA2(CSA2), .CSA1(CSA1), .CSA0(CSA0), .RSTA(RSTA),
    .CEB(CEB), .OCEB(OCEB), .CLKB(CLKB), .WEB(WEB), .CSB2(CSB2), .CSB1(CSB1), .CSB0(CSB0), .RSTB(RSTB)
);


DP16KD  #(
    .REGMODE_A("OUTREG"), .REGMODE_B("OUTREG")
) ebr_OUTREG_OUTREG (
    .DIA0(DIA[0]), .DIA1(DIA[1]), .DIA2(DIA[2]), .DIA3(DIA[3]), .DIA4(DIA[4]), .DIA5(DIA[5]), .DIA6(DIA[6]), .DIA7(DIA[7]), .DIA8(DIA[8]), .DIA9(DIA[9]), .DIA10(DIA[10]), .DIA11(DIA[11]), .DIA12(DIA[12]), .DIA13(DIA[13]), .DIA14(DIA[14]), .DIA15(DIA[15]), .DIA16(DIA[16]), .DIA17(DIA[17]),
    .DIB0(DIB[0]), .DIB1(DIB[1]), .DIB2(DIB[2]), .DIB3(DIB[3]), .DIB4(DIB[4]), .DIB5(DIB[5]), .DIB6(DIB[6]), .DIB7(DIB[7]), .DIB8(DIB[8]), .DIB9(DIB[9]), .DIB10(DIB[10]), .DIB11(DIB[11]), .DIB12(DIB[12]), .DIB13(DIB[13]), .DIB14(DIB[14]), .DIB15(DIB[15]), .DIB16(DIB[16]), .DIB17(DIB[17]),
    .ADA0(ADA[0]), .ADA1(ADA[1]), .ADA2(ADA[2]), .ADA3(ADA[3]), .ADA4(ADA[4]), .ADA5(ADA[5]), .ADA6(ADA[6]), .ADA7(ADA[7]), .ADA8(ADA[8]), .ADA9(ADA[9]), .ADA10(ADA[10]), .ADA11(ADA[11]), .ADA12(ADA[12]), .ADA13(ADA[13]),
    .ADB0(ADB[0]), .ADB1(ADB[1]), .ADB2(ADB[2]), .ADB3(ADB[3]), .ADB4(ADB[4]), .ADB5(ADB[5]), .ADB6(ADB[6]), .ADB7(ADB[7]), .ADB8(ADB[8]), .ADB9(ADB[9]), .ADB10(ADB[10]), .ADB11(ADB[11]), .ADB12(ADB[12]), .ADB13(ADB[13]),
    .DOA0(DOA_I[3][0]), .DOA1(DOA_I[3][1]), .DOA2(DOA_I[3][2]), .DOA3(DOA_I[3][3]), .DOA4(DOA_I[3][4]), .DOA5(DOA_I[3][5]), .DOA6(DOA_I[3][6]), .DOA7(DOA_I[3][7]), .DOA8(DOA_I[3][8]), .DOA9(DOA_I[3][9]), .DOA10(DOA_I[3][10]), .DOA11(DOA_I[3][11]), .DOA12(DOA_I[3][12]), .DOA13(DOA_I[3][13]), .DOA14(DOA_I[3][14]), .DOA15(DOA_I[3][15]), .DOA16(DOA_I[3][16]), .DOA17(DOA_I[3][17]),
    .DOB0(DOB_I[3][0]), .DOB1(DOB_I[3][1]), .DOB2(DOB_I[3][2]), .DOB3(DOB_I[3][3]), .DOB4(DOB_I[3][4]), .DOB5(DOB_I[3][5]), .DOB6(DOB_I[3][6]), .DOB7(DOB_I[3][7]), .DOB8(DOB_I[3][8]), .DOB9(DOB_I[3][9]), .DOB10(DOB_I[3][10]), .DOB11(DOB_I[3][11]), .DOB12(DOB_I[3][12]), .DOB13(DOB_I[3][13]), .DOB14(DOB_I[3][14]), .DOB15(DOB_I[3][15]), .DOB16(DOB_I[3][16]), .DOB17(DOB_I[3][17]),
    .CEA(CEA), .OCEA(OCEA), .CLKA(CLKA), .WEA(WEA), .CSA2(CSA2), .CSA1(CSA1), .CSA0(CSA0), .RSTA(RSTA),
    .CEB(CEB), .OCEB(OCEB), .CLKB(CLKB), .WEB(WEB), .CSB2(CSB2), .CSB1(CSB1), .CSB0(CSB0), .RSTB(RSTB)
);

assign DOA = DOA_I[sel];
assign DOB = DOB_I[sel];


endmodule