module vref (
  input in,
  output out
);

  assign out = in;

endmodule