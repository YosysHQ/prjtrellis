module top(input a, output q);
assign q = a;
endmodule
