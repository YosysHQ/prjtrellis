module top(output f);
    assign f = 1;
endmodule
