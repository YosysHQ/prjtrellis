module dcc_test1(input clki, input ce, output clko);

DCCA I1 (.CLKI (clki), .CE (ce), .CLKO (clko));

endmodule
