module top(
input TCK, TMS, TDI, JTDO2, JTDO1,
output TDO, JTDI, JTCK, JRTI2, JRTI1,
output JSHIFT, JUPDATE, JRSTN, JCE2, JCE1
);
    JTAGG jtag_i(.TCK(TCK), .TMS(TMS), .TDI(TDI), .JTDO2(JTDO2), .JTDO1(JTDO2),
       .TDO(TDO), .JTDI(JTDI), .JTCK(JTCK), .JRTI2(JRTI2), .JRTI1(JRTI1),
       .JSHIFT(JSHIFT), .JUPDATE(JUPDATE), .JRSTN(JRSTN), .JCE2(JCE2), .JCE1(JCE1));
endmodule
