module OB(input I, output O);
    assign O = I;
endmodule // OB
