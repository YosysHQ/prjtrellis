module OLVDS(input A, output Z, ZN);
    assign Z = A;
    assign ZN = ~A;
endmodule // OLVDS
