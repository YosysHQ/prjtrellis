module IB(input I, output O);
    assign O = I;
endmodule // IB
